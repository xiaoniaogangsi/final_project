module control_speed_motion