module Drawing_Engine(
//retrieve information from 