module frame_buffer ();


endmodule