module control_speed_motion();

endmodule
