module fire_control (input frame_Clk, Reset,
							input [7:0] keycode,
							output [9:0]  FireX, FireY);
							