module Drawing_Engine(